// adder_if.sv

interface adder_if;
 logic [1:0] a, b;
 logic cin;
 logic [1:0] sum;
 logic cout;
endinterface